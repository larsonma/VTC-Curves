*******************************************************
* Filename: RTL.cir
* Author: larsonma@msoe.edu <Mitchell Larson>
* Date: Apr 10 2018
* Provides:
* - DC analysis of a resistor-transistor logic circuit
* - originating in 1961
*******************************************************
.model npnt NPN BF=100 IS=1.8f


VA 1 0 DC 5
VCC 2 0 DC 5

RB 1 4 3.9K
RC 2 3 3.9K

Q1 3 4 0 npnt

.DC VA 0 5 0.001
.PROBE
.END

