*******************************************************
* Filename: CMOS.cir
* Author: larsonma@msoe.edu <Mitchell Larson>
* Date: Apr 10 2018
* Provides:
* - DC analysis of a MOSFET logic inverter circuit
* - originating in 1964
*******************************************************
.model pmod PMOS KP=80U VTO=-0.7V
.model nmod NMOS KP=200U VTO=0.6V

VA 1 0 DC 5
VDD 2 0 DC 5

M1 3 1 2 2 pmod W=10U L=2U
M2 3 1 0 0 nmod W=4U L=2U

.DC VA 0 5 0.001
.PROBE
.END

